*** SPICE deck for cell eor{sch} from library xyz
*** Created on Tue Apr 10, 2018 14:49:17
*** Last revised on Tue Apr 10, 2018 14:59:25
*** Written on Tue Apr 10, 2018 14:59:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 'D:\student\scmos18.mod'

.global gnd vdd

*** TOP LEVEL CELL: eor{sch}
Mnmos@2 s B net@64 gnd N L=0.4U W=0.4U
Mnmos@3 s nmos@3_g B gnd N L=0.4U W=0.4U
Mnmos@4 net@64 A gnd gnd N L=0.4U W=0.4U
Mpmos@2 A B s vdd P L=0.4U W=0.4U
Mpmos@3 B A s vdd P L=0.4U W=0.4U
Mpmos@4 vdd A net@64 vdd P L=0.4U W=0.4U


vdd vdd gnd 1.8v
vin A gnd pulse 0 1.8 0ns 1ps 1ps 1ns 2.002ns 50
vin1 B gnd pulse 0 1.8 0ns 1ps 1ps 2ns 4.002ns 50
.tran 0.02ns 50ns
.END
