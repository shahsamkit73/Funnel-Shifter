*** SPICE deck for cell mux{sch} from library xyz
*** Created on Sat Apr 07, 2018 12:38:34
*** Last revised on Tue Apr 10, 2018 15:35:38
*** Written on Tue Apr 10, 2018 15:35:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include 'D:\student\scmos18.mod'

.global gnd vdd

*** TOP LEVEL CELL: mux{sch}
Mnmos@11 A net@62 out gnd N L=0.4U W=0.4U
Mnmos@12 B S out gnd N L=0.4U W=0.4U
Mnmos@13 net@62 S gnd gnd N L=0.4U W=0.4U
Mpmos@11 out S A vdd P L=0.4U W=0.4U
Mpmos@12 out net@62 B vdd P L=0.4U W=0.4U
Mpmos@13 vdd S net@62 vdd P L=0.4U W=0.4U



vdd vdd gnd 1.8v
vin A gnd pulse 0 1.8 0ns 1ps 1ps 1ns 2.002ns 50
vin1 B gnd pulse 0 1.8 0ns 1ps 1ps 1ns 2.002ns 50
vin2 S gnd pulse 0 1.8 0ns 1ps 1ps 2ns 4.002ns 50
.tran 0.02ns 50ns
.END
